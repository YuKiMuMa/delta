library verilog;
use verilog.vl_types.all;
entity delta_vlg_vec_tst is
end delta_vlg_vec_tst;
